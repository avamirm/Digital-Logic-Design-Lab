module Adder(output[7:0] out,input[7:0]a);
	assign out = a + 8'd1;
endmodule
